library verilog;
use verilog.vl_types.all;
entity lab_1_2_vlg_vec_tst is
end lab_1_2_vlg_vec_tst;
