library verilog;
use verilog.vl_types.all;
entity lab_1_2_vlg_check_tst is
    port(
        UPS             : in     vl_logic;
        signal_sound    : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab_1_2_vlg_check_tst;
