module task1(

);

endmodule
